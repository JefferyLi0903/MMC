//`define SIM_PROFILE