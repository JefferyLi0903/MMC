//`define SIM_PROFILE
`define ethernet_IQ_output